library ieee;   --maiyyan saiyyan
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- ENABLES FOR PIPELINES
    
enTITy Controller is
    port(    
        CLK : in std_logic;
        Current_Zero, Current_Carry : in std_logic;
        New_Carry, New_Zero : in std_logic;
        IR : in std_logic_vector(15 downto 0); 
        Sign_Bit : in std_logic; -- hazard_beq signal -------- KARDE NA BHOSDIKE

        ZF_EN, CF_EN, RF_D3_EN, RF_PC_EN, SH_EN : out std_logic;
        MUX_SE_SEL, MUX_RF_D3_SEL, MUX_ALU1B_SEL, MUX_MEMDOUT_SEL, MUX_LM_SEL, MUX_DEST2_SEL, MUX_RF_A3_SEL : out std_logic;
        MUX_PC_SEL, MUX_DEST_SEL, MUX_ALU_A_SEL : out std_logic_vector(1 downto 0);
        MUX_ALU_B_SEL : out std_logic_vector(2 downto 0);
        ALU_OP :out std_logic_vector(3 downto 0)
    ); 
end enTITy;

architecture Struct of Controller is

type arr_2d is array (0 to 5, 15 downto 0) of std_logic;
signal Instructions : arr_2d : ("1011000000000000", "1011000000000000", "1011000000000000",
                       "1011000000000000", "1011000000000000", "1011000000000000");

signal IR_fetched : std_logic_vector(15 downto 0) : "1011000000000000";
shared variable prev3carry : std_logic_vector(0 to 2) := "000";
shared variable prev3zero : std_logic_vector(0 to 2) := "000";
shared variable is_lm, is_sm : std_logic_vector(1 downto 0) := "00";
shared variable shift_instr_en_lm : std_logic := '0';

begin 

IR_fetched <= IR;

process instruction_update(CLK)
begin
    if ( rising_edge(clk) ) then
        if(shift_instr_en_lm = '1') then
            Instructions(1 to 2) := Instructions(0 to 1);
            Instructions(0) := IR_fetched;
            Instructions(4 to 5) := Instructions(3 to 4);
        else 
            Instructions(1 to 5) := Instructions(0 to 4);
            Instructions(0) := IR_fetched;
        end if;
    else
        null;
    end if;
end process

process set_controls_stage1(CLK, Instructions, Sign_Bit)
begin
    if rising_edge(clk) then
        if ((Instructions(1, 15 downto 12) = "0110" or Instructions(1, 15 downto 12) = "0111" ) or is_lm(0) ) then --LM SM
            Instructions(0) := "1011000000000000";
            is_lm(0) := '1';
            RF_PC_EN <= '0';
        else
            is_lm(0) := '0';
            RF_PC_EN <= '1';
        end if;

 --     if (( Instructions(3, 15 downto 12) = "1000" or Instructions(3, 15 downto 12) = "1001" or Instructions(3, 15 downto 12) = "1010" ) and Sign_Bit = '1') or ( Instructions(3, 15 downto 12) = "1100") then -- BLT BLE BEQ or JAL
        if (( Instructions(3, 15 downto 12) = "1000" or Instructions(3, 15 downto 12) = "1001" or Instructions(3, 15 downto 12) = "1010" ) and Sign_Bit = '1')  then --changed for JAL
            MUX_PC_SEL <= "01";
            Instructions(0 to 2)="1011000000000000";
        elsif  ( Instructions(1, 15 downto 12) = "1100") then
            MUX_PC_SEL <= "01";
            Instruction(0)="1011000000000000";
        elsif Instructions(2, 15 downto 12) = "1101" then
            MUX_PC_SEL <= "10";
            Instructions(0 to 1)="1011000000000000";
        elsif Instructions(3, 15 downto 12) = "1111" then
            MUX_PC_SEL <= "11";
            Instructions(0 to 2)="1011000000000000";
        else 
            MUX_PC_SEL <= "00";
            -- LATCH
        end if;
    else
        null;
    end if; 
    
end process

process set_controls_stage2(CLK, Instructions)
begin
    if rising_edge(clk) then
        if ( is_sm = '1' ) then
            MUX_SM_SEL <= '1';
        else
            MUX_SM_SEL <= '0';
        end if;

        if ( Instructions(1, 15 downto 12) = "0011" or Instructions(1, 15 downto 12) = "0110" or Instructions(1, 15 downto 12) = "0111" or Instructions(1, 15 downto 12) = "1100" or Instructions(1, 15 downto 12) = "1111") then 
            MUX_SE_SEL <= "1";
        else 
            MUX_SE_SEL <= "0"; -- SE_6 IS DEFAULT
        end if;

        if ( Instructions(1, 15 downto 12) = "1000" or Instructions(1, 15 downto 12) = "1001" or Instructions(1, 15 downto 12) = "1010" or Instructions(1, 15 downto 12) = "1100" or Instructions(1, 15 downto 12) = "1111"  ) then 
           SH_EN <= "1";
        else      
           SH_EN <= "0";
        end if; 

    else
        null
    end if;
    
end process

process set_controls_stage3(CLK, Instructions)
begin

    variable opcode := Instructions(5, 15 downto 12)
    variable last3bits :=Instructions(5, 2 downto 0)

    if rising_edge(clk) then 
        if ( is_sm = '1' ) then --------------------------HAVE TO CHANGE 
            MUX_RF_A3_SEL <= '1';
        else
            MUX_RF_A3_SEL <= '0';
        end if;

        if (opcode = "0101" or opcode = "0111" or opcode = "1000" or opcode = "1111" or opcode = "1011") then -- SW, SM, BEQ, JRI or NOP then dont give enable
            RF_D3_EN <= "0"
        elsif ((opcode = "0001" and last3bits="010") or (opcode = "0001" and last3bits="110") or (opcode = "0010" and last3bits="010") or (opcode = "0010" and last3bits="110") ) and (prev3carry(2) = '0') -- ADC, ACC, NDC, NCC
            RF_D3_EN <= "0"
        elsif ((opcode = "0001" and last3bits="001") or (opcode = "0001" and last3bits="101") or (opcode = "0010" and last3bits="001") or (opcode = "0010" and last3bits="101") ) and (prev3zero(2) = '0') -- ADZ, ACZ, NDZ, NCZ
            RF_D3_EN <= "0";
        else
            RF_D3_EN <= "1";
        end if;

        if (opcode = "1100" or opcode = "1101") then -- JAL AND JLR
           MUX_RF_D3_SEL <= "1";
        else 
            MUX_RF_D3_SEL <= "0";
        end if;

        if (Instructions(2, 15 downto 12) = "0001" or Instructions(2, 15 downto 12) = "0010") then -- 5 to 3
            MUX_DEST_SEL <= "00";
        elsif (Instructions(2, 15 downto 12) = "0000" ) -- 8 to 6
            MUX_DEST_SEL <= "01";
        elsif (Instructions(2, 15 downto 12) = "0011" or Instructions(2, 15 downto 12) = "0100" or Instructions(2, 15 downto 12) = "1100" or Instructions(2, 15 downto 12) = "1101") -- 11 to 9
            MUX_DEST_SEL <= "10";
        else 
            null
        end if;

        if () then -- RA as it is
            MUX_ALU_A_SEL <= "00" 
        elsif () -- ALU1_C
            MUX_ALU_A_SEL <= "01"
        elsif () -- MEM_DOUT
            MUX_ALU_A_SEL <= "10"
        else -- WB_Forwarding
            MUX_ALU_A_SEL <= "11"
        end if;

        if () then -- Rb as it is
            MUX_ALU_B_SEL <= "000" 
        elsif () -- Normal IMM
            MUX_ALU_B_SEL <= "001"
        elsif () -- ALU_C
            MUX_ALU_B_SEL <= "010"
        elsif () -- MEM_DOUT
            MUX_ALU_B_SEL <= "011"
        else -- WB_Forwarding
            MUX_ALU_B_SEL <= "111"
        end if;

        if (is_lm(1) = '1') then -- Then LM has reached EX
            MUX_LM_SEL <= '1';
        else
            MUX_LM_SEL <= '0';
        end if;

    else 
        null
    end if;
end process

process set_controls_stage4(CLK, Instructions, Current_Carry, Current_Zero)
begin
    variable opcode := Instructions(3, 15 downto 12)
    variable last3bits :=Instructions(3, 2 downto 0)

    if ( Instructions(3, 15 downto 12) = "0110" ) then
        is_lm(1) := '1';
        shift_instr_enable := '1';
    else
        is_lm(1) := '0';
        shift_instr_enable := '0';
    end if;

    if (is_lm(1) = '1') then
        MUX_DEST2_SEL <= '1';
    else
        MUX_DEST2_SEL <= '0';
    end if;

    if (opcode="0001" and last3bits = "000") or (opcode = "0000") then 
        ZF_EN <= '1';
        CF_EN <= '1';
        ALU_OP <= "0000";
    elsif (opcode="0001" and last3bits = "010") then 
        if Current_Carry = '1' then
            ZF_EN <= '1';
            CF_EN <= '1';
            ALU_OP <= "0000";
        else
            ZF_EN <= '0';
            CF_EN <= '0';
            ALU_OP <= "1111";
        end if;
    elsif (opcode="0001" and last3bits = "001") then 
        if Current_Zero = '1' then
            ZF_EN <= '1';
            CF_EN <= '1';
            ALU_OP <= "0000";
        else
            ZF_EN <= '0';
            CF_EN <= '0';
            ALU_OP <= "1111";
        end if;
    elsif (opcode="0001" and last3bits = "011") then 
        ZF_EN <= '1';
        CF_EN <= '1';
        ALU_OP <= "0001";
    elsif (opcode="0001" and last3bits = "100") then 
        ZF_EN <= '1';
        CF_EN <= '1';
        ALU_OP <= "0010";
    elsif (opcode="0001" and last3bits = "110") then 
        if Current_Carry = '1' then
            ZF_EN <= '1';
            CF_EN <= '1';
            ALU_OP <= "0010";
        else
            ZF_EN <= '0';
            CF_EN <= '0';
            ALU_OP <= "1111";
        end if;
    elsif (opcode="0001" and last3bits = "101") then 
        if Current_Zero = '1' then
            ZF_EN <= '1';
            CF_EN <= '1';
            ALU_OP <= "0010";
        else
            ZF_EN <= '0';
            CF_EN <= '0';
            ALU_OP <= "1111";
        end if;
    elsif (opcode="0001" and last3bits = "111") then 
        ZF_EN <= '1';
        CF_EN <= '1';
        ALU_OP <= "0011";
    ---------------
    elsif (opcode="0010" and last3bits = "000") then 
        ZF_EN <= '1';
        CF_EN <= '1';
        ALU_OP <= "0100";
    elsif (opcode="0010" and last3bits = "010") then 
        if Current_Carry = '1' then
            ZF_EN <= '1';
            CF_EN <= '1';
            ALU_OP <= "0100";
        else
            ZF_EN <= '0';
            CF_EN <= '0';
            ALU_OP <= "1111";
        end if;
    elsif (opcode="0010" and last3bits = "001") then 
        if Current_Zero = '1' then
            ZF_EN <= '1';
            CF_EN <= '1';
            ALU_OP <= "0100";
        else
            ZF_EN <= '0';
            CF_EN <= '0';
            ALU_OP <= "1111";
        end if;
    ----------
    elsif (opcode="0010" and last3bits = "100") then 
        ZF_EN <= '1';
        CF_EN <= '1';
        ALU_OP <= "0101";
    elsif (opcode="0010" and last3bits = "110") then 
        if Current_Carry = '1' then
            ZF_EN <= '1';
            CF_EN <= '1';
            ALU_OP <= "0101";
        else
            ZF_EN <= '0';
            CF_EN <= '0';
            ALU_OP <= "1111";
        end if;
    elsif (opcode="0010" and last3bits = "101") then 
        if Current_Zero = '1' then
            ZF_EN <= '1';
            CF_EN <= '1';
            ALU_OP <= "0101";
        else
            ZF_EN <= '0';
            CF_EN <= '0';
            ALU_OP <= "1111";
        end if;    
    elsif (opcode="0011") then 
        ZF_EN <= '0';
        CF_EN <= '0';
        ALU_OP <= "0000"
    elsif (opcode="0100") then 
        ZF_EN <= '0';
        CF_EN <= '0';
        ALU_OP <= "0000";
    elsif (opcode="0101") then 
        ZF_EN <= '0'
        CF_EN <= '0'
        ALU_OP <= "0000"
    elsif (opcode="0110") then --LM
        ZF_EN <= '0';
        CF_EN <= '0';
        ALU_OP <= "0000";
    elsif (opcode="0111") then --SM
        ZF_EN <= '0';
        CF_EN <= '0';
        ALU_OP <= "0000";
    elsif (opcode="1000") then --BEQ
        ZF_EN <= '0';
        CF_EN <= '0';
        ALU_OP <= "0110";
    elsif (opcode="1001" and ) then --BLT
        ZF_EN <= '0';
        CF_EN <= '0';
        ALU_OP <= "0111";
    elsif (opcode="1010") then --BLE
        ZF_EN <= '0';
        CF_EN <= '0';
        ALU_OP <= "1000";
    elsif (opcode="1100") then --JAL
        ZF_EN <= '0';
        CF_EN <= '0';
        ALU_OP <= "1111";
    elsif (opcode="1101") then --JLR
        ZF_EN <= '0';
        CF_EN <= '0';
        ALU_OP <= "1111";
    elsif (opcode="1111") then --JRI
        ZF_EN <= '0';
        CF_EN <= '0';
        ALU_OP <= "0000";
    end if;
end process

process update_prevcarry(clk, New_Carry, New_Zero)
begin
    if(rising_edge(clk)) then
        prev3carry(1 to 2) := prev3carry(0 to 1)
        prev3carry(0) := New_Carry
        prev3zero(1 to 2) := prev3zero(0 to 1)
        prev3zero(0) := New_Zero
    else
        null
    end if;
end process;

process set_controls_stage5(CLK, Instructions)
begin
    if rising_edge(clk) then
        variable opcode := Instructions(4, 15 downto 12)

        if (opcode="0101") or (opcode = "0111") then  -- SM, SW
            MEM_WR_EN <= '1';
        else
            MEM_WR_EN <= '0';
        end if;
        
    else 
        null
    end if; 
end process


process set_controls_stage6(CLK, Instructions)
begin
    if rising_edge(clk) then
        variable opcode := Instructions(5, 15 downto 12)

        if (opcode="0100") or (opcode = "0110") then  -- LW, LM
            MUX_MEMDOUT_SEL <= '0'; -- MEM_DOUT
        else
            MUX_MEMDOUT_SEL <= '1'; -- ALU_C
        end if;

    else 
        null
    end if; 
end process

process hazard(CLK,Instructions)
begin  
    
end process;
end architecture;